/*************************************************************************
   > File Name: i2s_tx_10xe_tb_top.sv
   > Description: This file defines the AXI-Stream interface signals and associated clocking blocks for I2S transmitter functionality.
   > Author: Muhammad Junaid Ramzan
   > Modified: Muhammad Junaid Ramzan
   > Mail: muhammad.junaid@10xengineers.ai
   ---------------------------------------------------------------
   Copyright   (c)2024 10xEngineers
   ---------------------------------------------------------------
************************************************************************/

`include "i2s_tx_10xe_axi_stream_intf.sv"
`include "i2s_tx_10xe_axi4_lite_intf.sv"
`include "i2s_tx_10xe_dut_intf.sv"